module rambo

// adds two numbers of type T
pub fn add<T>(a1 T, a2 T) int {
	return a1 + a2
}