module rambo

// returns whatever `t` is passed in
pub fn identity<T>(t T) T {
	return t
}