module rambo

pub fn is_even(n int) bool {
	return n % 2 == 0
}
