module rambo

// always does logical and of two booleans
pub fn and(val1 bool, val2 bool) bool {
	return val1 && val2
}