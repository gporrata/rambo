module rambo

// returns true if `n` is even
pub fn is_even(n int) bool {
	return n % 2 == 0
}
