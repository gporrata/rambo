module rambo

pub fn is_positive(num int) bool {
	return num >= 0
}
