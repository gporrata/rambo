module rambo

pub fn inc<T>(t T) T {
	return t + 1
}