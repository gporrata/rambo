module rambo

// returns true if `num` is negative
pub fn is_negative(num int) bool {
	return num < 0
}
