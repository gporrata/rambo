module rambo

// note: will T always be boolean?
pub fn and(val1 bool, val2 bool) bool {
	return val1 && val2
}