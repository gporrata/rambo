module rambo

// increments `t` by 1
pub fn inc<T>(t T) T {
	return t + 1
}