module rambo

fn add<T>(val1 T, val2 T) T {
	return T + T
}

fn and<T>(val1 T, val2 T) T {
	return T && T
}