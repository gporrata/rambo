module rambo

pub fn identity<T>(t T) T {
	return t
}