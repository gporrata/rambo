module rambo

pub fn add<T>(a1 T, a2 T) int {
	return a1 + a2
}