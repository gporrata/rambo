module rambo

// todo: separate into files

//pub fn add<T>(val1 T, val2 T) T {
//	return T + T
//}

pub fn and<T>(val1 T, val2 T) T {
	return T && T
}