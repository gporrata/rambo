module rambo

pub fn is_negative(num int) bool { 
	return num < 0
}
