module rambo

fn and<T>(val1 T, val2 T) T {
	return T && T
}