module rambo

// returns true if `n` is odd
pub fn is_odd(n int) bool {
	return n % 2 == 1
}
