module rambo

pub fn is_odd(n int) bool {
	return n % 2 == 1
}
