module rambo

// returns true if `num` is positive
pub fn is_positive(num int) bool {
	return num >= 0
}
